module mag_comp_df(A_eq_B, A_gt_B, A_lt_B,
                   A,B);

output A_eq_B;
output A_gt_B;
output A_lt_B;
input [3:0] A, B;

wire not_B1, not_B0, not_

endmodule